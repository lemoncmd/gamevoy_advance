module main

import cpu as _ { Cpu }

fn main() {
	_ := Cpu.new()
	println('Hello World!')
}
